module in_out (input rst, input wire[4:0] in, output reg[31:0] out);
always @* begin
	case(in)
		//5'h00: out <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		5'h00: out <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
		5'h01: out <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
		5'h02: out <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;
		5'h03: out <= 32'b0000_0000_0000_0000_0000_0000_0000_1000; 
		5'h04: out <= 32'b0000_0000_0000_0000_0000_0000_0001_0000; 
		5'h05: out <= 32'b0000_0000_0000_0000_0000_0000_0010_0000; 
		5'h06: out <= 32'b0000_0000_0000_0000_0000_0000_0100_0000; 
		5'h07: out <= 32'b0000_0000_0000_0000_0000_0000_1000_0000; 
		5'h08: out <= 32'b0000_0000_0000_0000_0000_0001_0000_0000; 
		5'h09: out <= 32'b0000_0000_0000_0000_0000_0010_0000_0000; 
		5'h0A: out <= 32'b0000_0000_0000_0000_0000_0100_0000_0000; 
		5'h0B: out <= 32'b0000_0000_0000_0000_0000_1000_0000_0000; 
		5'h0C: out <= 32'b0000_0000_0000_0000_0001_0000_0000_0000; 
		5'h0D: out <= 32'b0000_0000_0000_0000_0010_0000_0000_0000; 
		5'h0E: out <= 32'b0000_0000_0000_0000_0100_0000_0000_0000; 
		5'h0F: out <= 32'b0000_0000_0000_0000_1000_0000_0000_0000; 
		5'h10: out <= 32'b0000_0000_0000_0001_0000_0000_0000_0000; 
		5'h11: out <= 32'b0000_0000_0000_0010_0000_0000_0000_0000; 
		5'h12: out <= 32'b0000_0000_0000_0100_0000_0000_0000_0000; 
		5'h13: out <= 32'b0000_0000_0000_1000_0000_0000_0000_0000; 
		5'h14: out <= 32'b0000_0000_0001_0000_0000_0000_0000_0000; 
		5'h15: out <= 32'b0000_0000_0010_0000_0000_0000_0000_0000; 
		5'h16: out <= 32'b0000_0000_0100_0000_0000_0000_0000_0000; 
		5'h17: out <= 32'b0000_0000_1000_0000_0000_0000_0000_0000; 
		5'h18: out <= 32'b0000_0001_0000_0000_0000_0000_0000_0000; 
		5'h19: out <= 32'b0000_0010_0000_0000_0000_0000_0000_0000; 
		5'h1A: out <= 32'b0000_0100_0000_0000_0000_0000_0000_0000; 
		5'h1B: out <= 32'b0000_1000_0000_0000_0000_0000_0000_0000; 
		5'h1C: out <= 32'b0001_0000_0000_0000_0000_0000_0000_0000; 
		5'h1D: out <= 32'b0010_0000_0000_0000_0000_0000_0000_0000; 
		5'h1E: out <= 32'b0100_0000_0000_0000_0000_0000_0000_0000; 
		5'h1F: out <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;	
		default: out<= 32'd123;
	endcase
	if (rst) begin
		out <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
	end
end 
endmodule 
